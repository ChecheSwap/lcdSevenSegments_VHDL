LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BASE IS PORT(
	XCLK : IN STD_LOGIC;
	XRST : IN STD_LOGIC;
	XRST2 : IN STD_LOGIC;
	
	XOUTPUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	XPOS: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);	
	XLED1 : OUT STD_LOGIC := '0';
	XLED2 : OUT STD_LOGIC := '0';
	XLED3 : OUT STD_LOGIC := '0';
	XLED4 : OUT STD_LOGIC := '0'
		
);
END BASE;

ARCHITECTURE BH OF BASE IS
	
	TYPE STATES IS (ZERO, ONE, TWO, THREE, FOUR , FIVE, SIX, SEVEN, EIGHT, NINE, STOP);
	SIGNAL STATE_NOW : STATES := ZERO;
	SIGNAL STATE_NEXT : STATES := ONE;
	
	CONSTANT SECOND : INTEGER := 1000000;	
	SIGNAL TIMESTAMP : INTEGER := SECOND;
	
	SIGNAL LEDSTATE : STD_LOGIC := '0';
	SIGNAL OUTPUT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');	
	

	CONSTANT BIN_ZERO : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000011";
	CONSTANT BIN_ONE : STD_LOGIC_VECTOR(7 DOWNTO 0) := "10011111";
	CONSTANT BIN_TWO : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00100101";
	CONSTANT BIN_THREE : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00001101";
	CONSTANT BIN_FOUR : STD_LOGIC_VECTOR(7 DOWNTO 0) := "10011001";
	CONSTANT BIN_FIVE : STD_LOGIC_VECTOR(7 DOWNTO 0) := "01001001";
	CONSTANT BIN_SIX : STD_LOGIC_VECTOR(7 DOWNTO 0) := "01000001";
	CONSTANT BIN_SEVEN : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011111";
	CONSTANT BIN_EIGHT : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000001";
	CONSTANT BIN_NINE : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00011001";	
	CONSTANT BIN_STOP : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";	
	
BEGIN
	
	BASE_TIME: PROCESS(XCLK, XRST, XRST2) 
	
		VARIABLE ENABLE_TIME : INTEGER := 0;	
		
		BEGIN		

			IF XRST = '0'  OR XRST2 = '0' THEN
				ENABLE_TIME := 0; 
				STATE_NOW <= STOP;	

			ELSIF  XCLK'EVENT AND XCLK = '1' THEN			
				IF(ENABLE_TIME >= TIMESTAMP) THEN
					ENABLE_TIME := 0;
					LEDSTATE <= NOT LEDSTATE;										
					STATE_NOW <= STATE_NEXT;														
				END IF;			

				ENABLE_TIME := ENABLE_TIME + 1;			
			END IF;

			IF XRST = '1' AND XRST2 = '1' THEN
				IF STATE_NOW = STOP THEN
					STATE_NOW <= ZERO;
				END IF;
			END IF;

	END PROCESS;
		
	
	ASS_NUMBER: PROCESS(XCLK, XRST, STATE_NOW) BEGIN
			
			CASE STATE_NOW IS
				WHEN ZERO => OUTPUT <= BIN_ZERO; 
				WHEN ONE => OUTPUT <= BIN_ONE;
				WHEN TWO => OUTPUT <= BIN_TWO;
				WHEN THREE => OUTPUT <= BIN_THREE;
				WHEN FOUR => OUTPUT <= BIN_FOUR;
				WHEN FIVE => OUTPUT <= BIN_FIVE;
				WHEN SIX => OUTPUT <= BIN_SIX;
				WHEN SEVEN => OUTPUT <= BIN_SEVEN;
				WHEN EIGHT => OUTPUT <= BIN_EIGHT;
				WHEN NINE => OUTPUT <= BIN_NINE;
				WHEN STOP => OUTPUT <= BIN_STOP;
			END CASE;
			
	END PROCESS;
	
	CALC_STATE : PROCESS(STATE_NOW) BEGIN
	
			CASE STATE_NOW IS				
				WHEN ZERO => STATE_NEXT <= ONE;
				WHEN ONE => STATE_NEXT <= TWO;
				WHEN TWO => STATE_NEXT <= THREE;
				WHEN THREE => STATE_NEXT <= FOUR;
				WHEN FOUR => STATE_NEXT <= FIVE;
				WHEN FIVE => STATE_NEXT <= SIX;
				WHEN SIX => STATE_NEXT <= SEVEN; 
				WHEN SEVEN => STATE_NEXT <= EIGHT;
				WHEN EIGHT => STATE_NEXT <= NINE;
				WHEN NINE => STATE_NEXT <= ZERO;
				WHEN OTHERS => STATE_NEXT <= ZERO;
			END CASE;
			
	END PROCESS;
	
	XLED1 <= LEDSTATE;
	XLED2 <= NOT LEDSTATE;
	XLED3 <= NOT LEDSTATE;
	XLED4 <= LEDSTATE;
	XOUTPUT <= OUTPUT;	
	XPOS <= "0000";
		
END BH;

 